`timescale 1ns / 1ps

module tb_int_to_fp;

    // 1. 信号定义
    reg         tb_clk;       // 用于控制测试流程的时钟
    reg  [63:0] tb_int_in;    // 输入：64位有符号整数
    wire [63:0] tb_fp_out;    // 输出：64位双精度浮点数

    // 2. 实例化待测模块 (DUT)
    // 根据你提供的接口定义，该模块为纯组合逻辑
    int_to_fp uut (
        .int_in     (tb_int_in),
        .fp_out     (tb_fp_out)
    );

    // 3. 时钟生成 (用于测试流程控制，非DUT必须)
    always #5 tb_clk = ~tb_clk;

    // 4. 定义测试任务
    task run_test;
        input [63:0] i_val;       // 输入整数
        input [63:0] expected;    // 预期浮点十六进制
        input [511:0] test_name;  // 测试名称
        
        begin
            // 建立输入
            tb_int_in = i_val;
            
            // 等待逻辑传播 (由于是组合逻辑，给一点延时即可，这里配合时钟边沿)
            @(posedge tb_clk);
            #1; //在此稍微延迟以确保信号稳定

            // 结果检查
            // 注意：浮点数比对通常不建议直接 ==，但对于整形转浮点，结果通常是确定的位模式
            if (tb_fp_out === expected) begin
                $display("PASS: %-45s. In=%d (0x%h) -> Got=0x%h", 
                         test_name, $signed(i_val), i_val, tb_fp_out);
            end else begin
                $display("FAIL: %-45s. In=0x%h, Expected=0x%h, Got=0x%h", 
                         test_name, i_val, expected, tb_fp_out);
            end
            
            // 插入间隙
            @(posedge tb_clk);
        end
    endtask

    // 5. 测试主流程
    initial begin
        // 初始化
        tb_clk = 0;
        tb_int_in = 0;

        // 生成波形文件
        $dumpfile("tb_int_to_fp.vcd");
        $dumpvars(0, tb_int_to_fp);

        #20;
        $display("================== 开始测试 int_to_fp ==================");
        $display("Rounding Mode: Round to Nearest, Ties to Even (Balanced)");

        // ------------------------------------------------------------
        // 组 1: 基础数值 (无需舍入)
        // ------------------------------------------------------------
        
        // Test 1: 0 -> 0.0
        run_test(64'd0, 64'h0000000000000000, 
                 "Test 1: Zero");

        // Test 2: 1 -> 1.0 (0x3FF0...0)
        run_test(64'd1, 64'h3FF0000000000000, 
                 "Test 2: Positive One");

        // Test 3: -1 -> -1.0 (0xBFF0...0)
        // -1 的补码是 0xFFFFFFFFFFFFFFFF
        run_test(-64'd1, 64'hBFF0000000000000, 
                 "Test 3: Negative One");

        // Test 4: 大的正数 (精确值)
        // 2^52 = 4,503,599,627,370,496 -> Exponent 1023+52, Mantissa 0
        run_test(64'h0010000000000000, 64'h4330000000000000, 
                 "Test 4: Large Exact Power of 2 (2^52)");

        // Test 5: 负的大数 (精确值)
        // -5 -> -5.0 (0xC014000000000000)
        run_test(-64'd5, 64'hC014000000000000, 
                 "Test 5: Small Negative Integer (-5)");

        // ------------------------------------------------------------
        // 组 2: 64位整数极值
        // ------------------------------------------------------------

        // Test 6: 最小负整数 (Min Int64)
        // -2^63 (0x8000...)。这是一个精确的2的幂次，可以精确表示。
        // Exp = 1023 + 63 = 1086 (0x43E). Sign = 1.
        run_test(64'h8000000000000000, 64'hC3E0000000000000, 
                 "Test 6: Int64 Min (-2^63)");

        // Test 7: 最大正整数 (Max Int64)
        // 2^63 - 1 (0x7FFF...). 双精度只有53位精度，需要舍入。
        // 值接近 2^63，且向偶数/最近舍入会进位变成 2^63。
        // 0x7FFF...FF -> 进位 -> 2^63 -> Exp 0x43E, Mantissa 0
        run_test(64'h7FFFFFFFFFFFFFFF, 64'h43E0000000000000, 
                 "Test 7: Int64 Max (Rounds up to 2^63)");

        // ------------------------------------------------------------
        // 组 3: 平衡舍入 (Round to Nearest Even) 关键测试
        // ------------------------------------------------------------
        // 双精度浮点数有53位有效数字(含隐含位)。
        // 当整数超过 2^53 时，LSB 开始无法表示，需要舍入。
        
        // Test 8: 舍入到最近的偶数 (向下去掉)
        // 输入: 2^53 + 1 = 9007199254740993 (0x20000000000001)
        // 此时精度位在 bit 1 (值为2)。bit 0 (值为1) 是"0.5 ULP"，正好在中间。
        // 前一位 (bit 1) 是 0 (偶数)。
        // 规则: Halfway case, round to even -> 向下舍入到 2^53
        // 预期: 2^53 (0x4340000000000000)
        run_test(64'h20000000000001, 64'h4340000000000000, 
                 "Test 8: Tie to Even (Round Down/Truncate)");

        // Test 9: 舍入到最近的偶数 (向上进位)
        // 输入: 2^53 + 3 = 9007199254740995 (0x20000000000003)
        // 位于 2^53+2 和 2^53+4 之间。
        // LSB权重是2。bit 0 (1) 是中间值。
        // 当前LSB (bit 1) 是 1 (奇数)。
        // 规则: Halfway case, round to even -> 向上进位到 2^53+4
        // 预期: 2^53 + 4. Exp=53. Mantissa LSB权重是2，所以Mantissa值为2。
        // Hex: 0x4340000000000002
        run_test(64'h20000000000003, 64'h4340000000000002, 
                 "Test 9: Tie to Even (Round Up/Increment)");

        // Test 10: 普通进位测试 (分数部分 > 0.5 ULP)
        // ------------------------------------------------------------
        // 输入数值: 2^54 + 3
        // Hex: 64'h0040000000000003
        // 二进制: ... 0001 (bit 54) ... 0000 0011 (bit 1,0)
        //
        // 【精度分析】
        // 1. 双精度浮点数只有 53 位精度 (1位隐含 + 52位显式)。
        // 2. 输入最高位 (MSB) 在 bit 54。
        // 3. 能够表示的最低有效位 (LSB) 位置 = 54 - 52 = 2。
        //    这意味着：权重为 2^2 (即 4) 的位是最后一位能保留的位。
        //    权重为 2^1 (2) 和 2^0 (1) 的位将被丢弃。
        //
        // 【舍入逻辑】
        // 丢弃部分数值 = 3 (二进制 11)。
        // 当前 LSB 的权重 = 4。半个 LSB (0.5 ULP) = 2。
        // 因为 3 > 2 (即 丢弃值 > 0.5 ULP)，必须向上进位 (Round Up)。
        //
        // 【预期结果】
        // 目标值 = (2^54 + 3) 向上舍入到最近的 4 的倍数 => 2^54 + 4。
        // 2^54 + 4 的浮点表示：
        // 科学计数法: 1.00...001 * 2^54  (尾数最低位对应 4/2^54)
        // 指数 (Exp): 1023 + 54 = 1077 = 0x435
        // 尾数 (Mant): 最低位为1，其余为0 (即 52'h0000000000001)
        // 组合 Hex: 0x4350000000000001
        run_test(64'h0040000000000003, 64'h4350000000000001, 
                "Test 10: Round Up (Fraction > 0.5)");

        $display("================== 结束测试 int_to_fp ==================");
        #20;
        $finish;
    end

endmodule
